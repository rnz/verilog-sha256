/*****************************************************************************/
/*   SHA 256 module testbench, 512bit version                                */ 
/*   Aishwarya Nagarajan, UW-Madison, ERCBench Researcher                    */
/*   Inputs: clk, rst, valid,last, first, msg_in (512bits)                   */
/*   Outputs: ready, msg_out (256 bits)                                      */
/*****************************************************************************/

module t_sha_multi_chunks2();
   
   //declairng input and output regs and wires	   
   reg clk, rst, valid, first, last;
   reg [511:0] msg_in;
   wire [255:0] msg_out; 
   wire ready;
   
   //instatiating UUT	 
   sha_multi_chunks2 UUT (clk, rst,valid,first,last, msg_in, msg_out, ready);
   
   //creating clock
   initial clk=1'b0;
   always @(clk) clk<= #5 ~clk;
   
   //assigning inputs 
   initial begin
       rst = 1'b1; 
       valid = 1'b0;
       #11 rst = 1'b0;
       #10 valid = 1'b1;
       first = 1'b1;
       last = 1'b0; 
       msg_in = 512'b01100001_01100010_01100011_01100100_01100010_01100011_01100100_01100101_01100011_01100100_01100101_01100110_01100100_01100101_01100110_01100111_01100101_01100110_01100111_01101000_01100110_01100111_01101000_01101001_01100111_01101000_01101001_01101010_01101000_01101001_01101010_01101011_01101001_01101010_01101011_01101100_01101010_01101011_01101100_01101101_01101011_01101100_01101101_01101110_01101100_01101101_01101110_01101111_01101101_01101110_01101111_01110000_01101110_01101111_01110000_01110001_10000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
       #640 first = 1'b0;
       #5 last = 1'b1; 
       msg_in = 512'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_11000000; 
       #640 first = 1'b0;
       #5 last = 1'b1; 
       msg_in = 512'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_11000000; 
       #640 first = 1'b0;
       #5 last = 1'b1; 
       msg_in = 512'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_11000000; 
       #640 first = 1'b0;
       #5 last = 1'b1; 
       msg_in = 512'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_11000000; 
       #640 first = 1'b0;
       #5 last = 1'b1; 
       msg_in = 512'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_11000000; 
   end  

   //force simulation end
   initial begin
       #15000 $stop; 
   end
   
endmodule




